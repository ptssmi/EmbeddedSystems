`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/14/2020 09:53:42 PM
// Design Name: 
// Module Name: Main_TestBench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Main_TestBench(

    );
    


    
    reg [3:0] IN1;
    reg [3:0] IN2;
    wire  [3:0] OUT;
    wire  CF;
    wire  Z;
    reg [1:0] CTRL;
    reg CLK;
    
    
    
    
    
endmodule
